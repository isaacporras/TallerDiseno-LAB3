//MAIN
