module flag_negativo #(parameter N = 8)(
							input logic [N-1:0] ultimo_bit,
							output logic [N-1:0] resultado );
										
assign resultado = ultimo_bit;

endmodule 