module correr_derecha #(parameter N = 8)(input logic [N-1:0] A,
													  input logic [N-1:0] B,
													  output logic [N-1:0] shift_right_out);

assign shift_right_out = A >> B;


endmodule 